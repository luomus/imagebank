title = Bildbanken - Identifiera Finlands Arter | Finlands Artdatacenter