imagebank = Bildbanken
tagline = Identifiera Finlands Arter
finbif = Finlands Artdatacenter
finbif_short = FinBIF

documentation =  Instruktioner
support = Support och feedback
change_language = Change language | Byt språk

login = Logga in
logout =  Logga ut
logged_in_as = Inloggad som

menu_home = Startsida
menu_browse = Bläddra
menu_curate = Kvalitetskontroll
menu_admin = Admin
menu_taxon_select = Taxonval

error_header = Tyvärr! Något gick fel...

admin_main = Admin | Bildhantering
admin_single_title = Redigera en bild
admin_single_body = Ange bildens adress (t.ex. https://image.laji.fi/MM.123/kuva.jpg) eller bildens identifierare (t.ex. MM.123 eller http://tun.fi/MM.123)
admin_taxon_title = Redigera taxonbilder
admin_taxon_body = Ange taxonens identifierare (t.ex. MX.123) eller dess vetenskapliga eller svenska namn
admin_select_image = Välj en bild att redigera
admin_info = <p>Admin-sektionen är ett underhållsverktyg och är inte avsett för vanlig artbildskuratering.</p><p>Här kan du redigera alla bilder, inklusive provbilder som lagts till i Kotka och observationsbilder som lagts till via Vihko.</p><p>Du kan redigera alla bildinformationer som inte kan ändras i artbildssektionen, t.ex. licens, fotografens namn och nyckelord.</p><p>Du kan även helt ta bort bilder.</p><p>I fall av avsiktlig missbruk eller skadegörelse, är det bättre att annotera observationen med en Spam-tag.</p>

taxon_autocomplete_placeholder = Par apollo, L dryas, Metalimnobia, knölsvan, MX.123
select_taxon = Välj taxon
exact_matches = Exakta träffar
partial_matches = Partiella träffar
likely_matches = Troliga träffar
no_taxon_matches = Inga träffar för sökordet
taxon_search_term = Matchar med sökterm
no_images = Inga bilder
edit_image = Redigera bild

must_be_admin = Du är inte inloggad eller saknar behörighet!
unknown_taxon = Okänd taxon-ID!
unknown_image = Okänd media-ID!