imagebank = Bildbanken
tagline = Identifiera Finlands Arter
finbif = Finlands Artdatacenter
finbif_short = FinBIF

documentation =  Instruktioner
support = Support och feedback

login = Logga in
logout =  Logga ut

menu_browse = Bläddra
menu_curate = Kvalitetskontroll
menu_admin = ADMIN
