imagebank = Bildbanken
tagline = Identifiera Finlands Arter
finbif = Finlands Artdatacenter
finbif_short = FinBIF

documentation =  Instruktioner
support = Support och feedback
change_language = Change language | Byt språk

login = Logga in
logout =  Logga ut
logged_in_as = Inloggad som

menu_home = Startsida
menu_browse = Bläddra
menu_curate = Kvalitetskontroll
menu_admin = Admin
menu_taxon_select = Taxonval

error_header = Tyvärr! Något gick fel...

admin_main = Admin | Bildhantering
admin_single_title = Redigera en bild
admin_single_body = Ange bildens adress (t.ex. https://image.laji.fi/MM.123/kuva.jpg) eller bildens identifierare (t.ex. MM.123 eller http://tun.fi/MM.123)
admin_taxon_title = Redigera taxonbilder
admin_taxon_body = Ange taxonens identifierare (t.ex. MX.123) eller dess vetenskapliga eller svenska namn
admin_select_image = Välj en bild att redigera
admin_info = <p>Admin-sektionen är ett underhållsverktyg och är inte avsett för vanlig artbildskuratering.</p><p>Här kan du redigera alla bilder, inklusive provbilder som lagts till i Kotka och observationsbilder som lagts till via Vihko.</p><p>Du kan redigera alla bildinformationer som inte kan ändras i artbildssektionen, t.ex. licens, fotografens namn och nyckelord.</p><p>Du kan även helt ta bort bilder.</p>
admin_edit_image = Redigera bild
admin_delete_image = Ta bort bild
admin_delete_image_note = <p>Observera att om du tar bort en bild från ett prov/exemplar (Kotka, Vihko, Löydös), kommer observationen att behålla en "trasig bild".</p><p>För Kotka provbilder kommer borttagningen av bilden att fördröjas i sökresultaten tills proverna omindexeras.</p><p>Bildborttagning skickas inte till Laji.fi datalagret, så där kommer den trasiga bilden att finnas kvar tills observationen redigeras.</p><p>För artbilder kan bilden ha valts för Pinkka, och där visas den trasiga bilden.</p><p>Det säkraste sättet att ta bort en artbild är att lämna bilden intakt och ta bort taksonidentifieraren/identifierarna från den.</p><p>I fall av avsiktlig missbruk eller skadegörelse, är det bättre att annotera observationen med en Spam-tag.</p>
admin_delete_confirm = Är du säker på att du vill ta bort denna bild?

taxon_autocomplete_placeholder = Par apollo, L dryas, Metalimnobia, knölsvan, MX.123
select_taxon = Välj taxon
exact_matches = Exakta träffar
partial_matches = Partiella träffar
likely_matches = Troliga träffar
no_taxon_matches = Inga träffar för sökordet
taxon_search_term = Matchar med sökterm

no_images = Inga bilder

save = Spara
save_success = Sparat!
cancel = Ångra
cancel_confirm = Är du säker på att du vill ångra alla ändringar?

yes = Ja
no = Nej

must_be_admin = Du är inte inloggad eller saknar behörighet!
unknown_taxon = Okänd taxon-ID!
unknown_image = Okänd media-ID!

group_authors = Författare
label_capturers = Fotograf
label_rightsOwner = Licensägare
label_license = Licens

group_dates = Datum
label_captureDateTime = Registreringstidpunkt
label_uploadDateTime = Uppladdningstidpunkt

group_taxon_images = Taxonbilder
label_taxonIds = Taxon-ID
label_verbatim = Verbatim
label_primaryForTaxon = Primär för taxon
label_type = Typ
label_sex = Kön
label_lifeStage = Livsfas
label_plantLifeStage = Växtens livsfas
label_side = Sida

group_captions = Bildtexter
label_caption = Bildtext
label_taxonDescriptionCaptionFI = Taxonbeskrivningstext - FI
label_taxonDescriptionCaptionSV = Taxonbeskrivningstext - SV
label_taxonDescriptionCaptionEN = Taxonbeskrivningstext - EN

group_misc = Övrigt
label_documentIds = Dokument-ID
label_tags = Nyckelord
label_sortOrder = Sorteringsordning

group_unmodifiable = Oföränderliga fält
label_sourceSystem = Källsystem
label_uploadedBy = Uppladdad av
label_secret = Hemlig
label_originalFilename = Ursprungligt filnamn
label_fullResolutionMediaAvailable = Fullupplöst media tillgänglig (via dataförfrågan)
