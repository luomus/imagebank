imagebank = Bildbanken
tagline = Identifiera Finlands Arter
finbif = Finlands Artdatacenter
finbif_short = FinBIF
privacy_policy = Integritetspolicy
privacy_policy_link = https://laji.fi/privacypolicy
accessibility_statement = NOP
accessibility_statement_link = NOP
finbif_mission = Finlands Artdatacenter samlar och förenar finländska artinformationsdata som en konsekvent och öppen enhet för forskning och utbildning, förvaltning och den breda allmänheten.

documentation =  Instruktioner
doc_link = https://info.laji.fi/en/frontpage/instructions-to-species-image-management-image-bank/
support = Support och feedback
change_language = Change language | Byt språk

login = Logga in
logout =  Logga ut
logged_in_as = Inloggad som

menu_home = Startsida
menu_browse = Bläddra
menu_curate = Kvalitetskontroll
menu_admin = Admin
menu_taxon_select = Taxonval
menu_image_select = Bildval

error_header = Tyvärr! Något gick fel...

browse_title = Bläddra | Bläddring och innehållsskapande
curate_title = Kvalitetskontroll | Bildkuratering

preferences = Inställningar
group = Organismgrupp
group_select = Välj en organismgrupp  
order = Ordning
taxonomic = Taxonomisk
alphabetic = Alfabetisk
taxa_preference = Finska arter 
taxa_finnish = Endast finska
taxa_all = Alla
taxon_ranks_preference = Taxonomiska nivåer
category_filter = Kategorier
uncategorized = Okategoriserad
page_size = Sidstorlek
image_size = Bildstorlek
image_size_small = Liten
image_size_large = Stor
content_creation_preference = Innehållsskapande
on = På
off = Av
close = Stäng
open = Öppna
no_matches = Inga resultat matchar
show_more = Visa mer
change = Ändra
select = Välj
edit = Redigera

taxon_tree = Taxonomiska nivåer
taxon_tree_no_taxa = Inga taxon att visa på denna nivå

admin_main = Admin | Bildhantering
admin_single_title = Redigera en bild
admin_single_body = Ange bildens adress (t.ex. https://image.laji.fi/MM.123/kuva.jpg) eller bildens identifierare (t.ex. MM.123 eller http://tun.fi/MM.123)
admin_taxon_title = Redigera taxonbilder
admin_taxon_body = Ange taxonens identifierare (t.ex. MX.123) eller dess vetenskapliga eller svenska namn
admin_add_image_title = Ladda upp bild
admin_add_image_title_multi = Ladda upp bilder
admin_add_image_info = Gå till taxonsidan för att lägga till flera bilder.
admin_select_image = Välj en bild att redigera
admin_info = <p>Admin-sektionen är ett underhållsverktyg och är inte avsett för vanlig artbildskuratering.</p><p>Här kan du redigera alla bilder, inklusive provbilder som lagts till i Kotka och observationsbilder som lagts till via Vihko.</p><p>Du kan redigera alla bildinformationer som inte kan ändras i artbildssektionen, t.ex. licens, fotografens namn och nyckelord.</p><p>Du kan även helt ta bort bilder.</p>
admin_edit_image = Redigera bild
admin_delete_image = Ta bort bild
admin_delete_image_note = <h5>Observera följande om borttagning av bilder:</h5><ul><li>Om du tar bort en prov- eller observationsbild (från Kotka, Vihko eller Löydös), lämnas en trasig bild kvar i observationen.</li><li>För Kotkas provbilder syns borttagningen inte omedelbart i sökresultaten, utan först när proverna har indexerats på nytt.</li><li>Information om borttagning av bilden överförs inte till Laji.fi-datalagret. Därför visas den trasiga bilden där tills observationen redigeras.</li><li>För artbilder kan bilden vara vald till Pinkka, och då visas den trasiga bilden även där.</li><li>I stället för att ta bort en artbild är det oftast säkrast att låta bilden vara kvar och i stället ta bort dess taxonidentifiering(ar).</li><li>Vid misstanke om vandalism räcker det inte att bara ta bort bilden. Markera dessutom observationen med Spam.</li></ul>
admin_delete_confirm = Är du säker på att du vill ta bort denna bild?
admin_delete_success = Borttagen!
admin_make_primary = Gör till primär för denna taxon
admin_tag_images = Tagga bilder
admin_tag_done = Klar/Uppdatera
admin_click_to_add_tags = Klicka på bilden för att lägga till taggar
admin_secret_image_help = En hemlig bild är inte offentligt tillgänglig. För att visa den krävs en speciell hemlig nyckel. Markera inte detta om du inte vet exakt varför.
admin_image_add_success = Uppladdad! Vänligen fyll i metadata såsom fotografens namn och licens.

taxon_autocomplete_placeholder = Par apollo, L dryas, Metalimnobia, knölsvan, MX.123
select_taxon = Välj taxon
exact_matches = Exakta träffar
partial_matches = Partiella träffar
likely_matches = Troliga träffar
no_taxon_matches = Inga träffar för sökordet
taxon_search_term = Matchar med sökterm

no_images = Inga bilder
no_image = Ingen bild
drop_image = Dra och släpp en bild här, eller klicka för att välja en.
drop_image_multi = Dra och släpp bilder här, eller klicka för att välja flera.

save = Spara
save_success = Sparat!
cancel = Ångra
cancel_confirm = Är du säker på att du vill ångra alla ändringar?
clear_all = Rensa alla

yes = Ja
no = Nej

loading = Belastning
esc_closes = stänger galleriet

must_be_admin = Du är inte inloggad eller saknar behörighet!
unknown_taxon = Okänd taxon-ID!
unknown_image = Okänd media-ID!
invalid_integer = Ogiltigt heltal
invalid_datetime = Ogiltigt datum/tidsformat
invalid_boolean = Ogiltigt värde, ska vara true/false
file_missing = Fil saknas!
file_too_large = Filen är för stor. Den maximala storleken är 50 MB.
invalid_parameters = Ogiltiga parametrar

group_authors = Författare
label_capturer = Fotograf
label_capturers = Fotografer
label_rightsOwner = Rättighetsinnehavare
label_license = Licens
label_captureDateTime = Registreringstidpunkt

group_taxon_images = Taxonbilder
label_taxonIds = Taxon-ID
label_verbatim = Verbatim
label_primaryForTaxon = Primär för taxon
label_type = Typ
label_sex = Kön
label_lifeStage = Livsfas
label_plantLifeStage = Växtens livsfas
label_side = Sida

group_captions = Bildtexter
label_caption = Bildtext
label_taxonDescriptionCaptionFI = Taxonbeskrivningstext - FI
label_taxonDescriptionCaptionSV = Taxonbeskrivningstext - SV
label_taxonDescriptionCaptionEN = Taxonbeskrivningstext - EN

group_misc = Övrigt
label_sortOrder = Sorteringsordning
sort_order_info = 0 = visas först, stora nummer visas senare
label_documentIds = Dokument-ID
label_tags = Nyckelord
label_fullResolutionMediaAvailable = Formulär för begäran om fullversion

group_unmodifiable = Oföränderliga fält
label_sourceSystem = Källsystem
label_uploadedBy = Uppladdad av
label_uploadDateTime = Uppladdningstidpunkt
label_modifiedBy = Ändrad av  
label_modifiedDateTime = Ändringstidpunkt
label_secret = Hemlig
label_originalFilename = Ursprungligt filnamn
